`ifndef DEFS
`define DEFS

`define MANUAL_DEBUG

`define UNIT_BCD_W      6
`define PULSE_CNT_W     40

`define MAX_MORSE_LEN   5
`define MORSE_LEN_W     3
`define CHAR_W          6
`define MAX_CHARS       6


`define CHAR_CODE_SPACE   `CHAR_W'd31

`define CHAR_CODE_0   `CHAR_W'd0
`define CHAR_CODE_1   `CHAR_W'd1
`define CHAR_CODE_2   `CHAR_W'd2
`define CHAR_CODE_3   `CHAR_W'd3
`define CHAR_CODE_4   `CHAR_W'd4
`define CHAR_CODE_5   `CHAR_W'd5
`define CHAR_CODE_6   `CHAR_W'd6
`define CHAR_CODE_7   `CHAR_W'd7
`define CHAR_CODE_8   `CHAR_W'd8
`define CHAR_CODE_9   `CHAR_W'd9
`define CHAR_CODE_A   `CHAR_W'd10
`define CHAR_CODE_B   `CHAR_W'd11
`define CHAR_CODE_C   `CHAR_W'd12
`define CHAR_CODE_D   `CHAR_W'd13
`define CHAR_CODE_E   `CHAR_W'd14
`define CHAR_CODE_F   `CHAR_W'd15


`define CHAR_ASCI_ARRAY  "0123456789ABCDEF                "

`define CHAR_MORSE_A   ".-"
`define CHAR_MORSE_B   "-..."
`define CHAR_MORSE_C   "-.-."
`define CHAR_MORSE_D   "-.."
`define CHAR_MORSE_E   "."
`define CHAR_MORSE_F   "..-."




`endif